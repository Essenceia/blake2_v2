module emulator(
	input wire clk, 
	output wire [7:0] segA_o
);

assign segA_o = 8'hFF;

endmodule
